//APB inerface 
